
module mem #(                   // 
    parameter  ADDR_LEN  = 11   // 
) (
    input  clk, rst,
    input  [ADDR_LEN-1:0] addr, // memory address
    output reg [31:0] rd_data,  // data read out
    input  wr_req,
    input  [31:0] wr_data       // data write in
);
localparam MEM_SIZE = 1<<ADDR_LEN;
reg [31:0] ram_cell [MEM_SIZE];

always @ (posedge clk or posedge rst)
    if(rst)
        rd_data <= 0;
    else
        rd_data <= ram_cell[addr];

always @ (posedge clk)
    if(wr_req) 
        ram_cell[addr] <= wr_data;

initial begin
    // dst matrix C
    ram_cell[       0] = 32'h0;  // 32'h529d69cb;
    ram_cell[       1] = 32'h0;  // 32'h02f94a71;
    ram_cell[       2] = 32'h0;  // 32'hbade3799;
    ram_cell[       3] = 32'h0;  // 32'hbb1c8c96;
    ram_cell[       4] = 32'h0;  // 32'hcb3a0b07;
    ram_cell[       5] = 32'h0;  // 32'h976ce6eb;
    ram_cell[       6] = 32'h0;  // 32'hcac30239;
    ram_cell[       7] = 32'h0;  // 32'h39a5f666;
    ram_cell[       8] = 32'h0;  // 32'haee5f5c5;
    ram_cell[       9] = 32'h0;  // 32'hdf7f4f64;
    ram_cell[      10] = 32'h0;  // 32'h705dcb87;
    ram_cell[      11] = 32'h0;  // 32'hc026e3b8;
    ram_cell[      12] = 32'h0;  // 32'h353a8c7d;
    ram_cell[      13] = 32'h0;  // 32'hc9624f4b;
    ram_cell[      14] = 32'h0;  // 32'hacaef33e;
    ram_cell[      15] = 32'h0;  // 32'h086b3ce3;
    ram_cell[      16] = 32'h0;  // 32'h825894ae;
    ram_cell[      17] = 32'h0;  // 32'h050c768f;
    ram_cell[      18] = 32'h0;  // 32'h329b1268;
    ram_cell[      19] = 32'h0;  // 32'h071f4c3f;
    ram_cell[      20] = 32'h0;  // 32'h0593157b;
    ram_cell[      21] = 32'h0;  // 32'hb9c72f6b;
    ram_cell[      22] = 32'h0;  // 32'h0f1f2d0f;
    ram_cell[      23] = 32'h0;  // 32'he07ef731;
    ram_cell[      24] = 32'h0;  // 32'hf49a40bd;
    ram_cell[      25] = 32'h0;  // 32'he2072d89;
    ram_cell[      26] = 32'h0;  // 32'h6c274d74;
    ram_cell[      27] = 32'h0;  // 32'h13aa2d00;
    ram_cell[      28] = 32'h0;  // 32'h71476c9f;
    ram_cell[      29] = 32'h0;  // 32'hf89df322;
    ram_cell[      30] = 32'h0;  // 32'h49019878;
    ram_cell[      31] = 32'h0;  // 32'h821fcab7;
    ram_cell[      32] = 32'h0;  // 32'hd5aa61b0;
    ram_cell[      33] = 32'h0;  // 32'h1638661b;
    ram_cell[      34] = 32'h0;  // 32'h7875ed22;
    ram_cell[      35] = 32'h0;  // 32'h3fae2d60;
    ram_cell[      36] = 32'h0;  // 32'h92bf4194;
    ram_cell[      37] = 32'h0;  // 32'ha52ad06e;
    ram_cell[      38] = 32'h0;  // 32'hcfa05581;
    ram_cell[      39] = 32'h0;  // 32'h4fa3c9fd;
    ram_cell[      40] = 32'h0;  // 32'h151c7172;
    ram_cell[      41] = 32'h0;  // 32'hcf53a99b;
    ram_cell[      42] = 32'h0;  // 32'hd6971e1b;
    ram_cell[      43] = 32'h0;  // 32'h3c8af1c4;
    ram_cell[      44] = 32'h0;  // 32'hd8c51060;
    ram_cell[      45] = 32'h0;  // 32'hc562e79d;
    ram_cell[      46] = 32'h0;  // 32'h33721152;
    ram_cell[      47] = 32'h0;  // 32'h818c6345;
    ram_cell[      48] = 32'h0;  // 32'h2e7ba987;
    ram_cell[      49] = 32'h0;  // 32'h71bd3114;
    ram_cell[      50] = 32'h0;  // 32'h0da02ecd;
    ram_cell[      51] = 32'h0;  // 32'hc4d8e1e9;
    ram_cell[      52] = 32'h0;  // 32'h49f021ba;
    ram_cell[      53] = 32'h0;  // 32'h0ec3b631;
    ram_cell[      54] = 32'h0;  // 32'hd4c2b7f4;
    ram_cell[      55] = 32'h0;  // 32'hc2b1225f;
    ram_cell[      56] = 32'h0;  // 32'hd31ce741;
    ram_cell[      57] = 32'h0;  // 32'habab1f29;
    ram_cell[      58] = 32'h0;  // 32'hcb24e9ce;
    ram_cell[      59] = 32'h0;  // 32'hdd02bfd1;
    ram_cell[      60] = 32'h0;  // 32'hec5a598a;
    ram_cell[      61] = 32'h0;  // 32'h94b493a5;
    ram_cell[      62] = 32'h0;  // 32'hf1f6ecf6;
    ram_cell[      63] = 32'h0;  // 32'h0a79ab5e;
    ram_cell[      64] = 32'h0;  // 32'h15f977d9;
    ram_cell[      65] = 32'h0;  // 32'h4e4a543b;
    ram_cell[      66] = 32'h0;  // 32'h982b68c3;
    ram_cell[      67] = 32'h0;  // 32'h7ac1bb7e;
    ram_cell[      68] = 32'h0;  // 32'hdc757760;
    ram_cell[      69] = 32'h0;  // 32'h2854a2a3;
    ram_cell[      70] = 32'h0;  // 32'h0fcc9b7b;
    ram_cell[      71] = 32'h0;  // 32'h09f90cf0;
    ram_cell[      72] = 32'h0;  // 32'hf25762e6;
    ram_cell[      73] = 32'h0;  // 32'h87f71e6b;
    ram_cell[      74] = 32'h0;  // 32'h7266c80d;
    ram_cell[      75] = 32'h0;  // 32'hd4ade938;
    ram_cell[      76] = 32'h0;  // 32'h633fb0d1;
    ram_cell[      77] = 32'h0;  // 32'h9defcd43;
    ram_cell[      78] = 32'h0;  // 32'hd08cdfc2;
    ram_cell[      79] = 32'h0;  // 32'hbdc75e41;
    ram_cell[      80] = 32'h0;  // 32'h30813e29;
    ram_cell[      81] = 32'h0;  // 32'ha0049212;
    ram_cell[      82] = 32'h0;  // 32'h06884a07;
    ram_cell[      83] = 32'h0;  // 32'h06255523;
    ram_cell[      84] = 32'h0;  // 32'heed3c6ef;
    ram_cell[      85] = 32'h0;  // 32'hefbea70a;
    ram_cell[      86] = 32'h0;  // 32'ha6ca84c7;
    ram_cell[      87] = 32'h0;  // 32'hb1ef6593;
    ram_cell[      88] = 32'h0;  // 32'ha6e9c962;
    ram_cell[      89] = 32'h0;  // 32'h2e78b11f;
    ram_cell[      90] = 32'h0;  // 32'h70f4ddc3;
    ram_cell[      91] = 32'h0;  // 32'hb8ba3756;
    ram_cell[      92] = 32'h0;  // 32'ha07bf12f;
    ram_cell[      93] = 32'h0;  // 32'he7abd703;
    ram_cell[      94] = 32'h0;  // 32'hf987f1d0;
    ram_cell[      95] = 32'h0;  // 32'h23e0b4bf;
    ram_cell[      96] = 32'h0;  // 32'h6f514a80;
    ram_cell[      97] = 32'h0;  // 32'h99d620da;
    ram_cell[      98] = 32'h0;  // 32'he4f84c99;
    ram_cell[      99] = 32'h0;  // 32'hb3a6ae46;
    ram_cell[     100] = 32'h0;  // 32'h8f61030a;
    ram_cell[     101] = 32'h0;  // 32'h68886d50;
    ram_cell[     102] = 32'h0;  // 32'h12df5208;
    ram_cell[     103] = 32'h0;  // 32'h86f8d7c8;
    ram_cell[     104] = 32'h0;  // 32'h16151bc1;
    ram_cell[     105] = 32'h0;  // 32'h84e78bab;
    ram_cell[     106] = 32'h0;  // 32'hb5ebdc3c;
    ram_cell[     107] = 32'h0;  // 32'h2027fc59;
    ram_cell[     108] = 32'h0;  // 32'hca1cd67c;
    ram_cell[     109] = 32'h0;  // 32'h1f464bf4;
    ram_cell[     110] = 32'h0;  // 32'hd3a26c4a;
    ram_cell[     111] = 32'h0;  // 32'h7a136e6a;
    ram_cell[     112] = 32'h0;  // 32'ha7610658;
    ram_cell[     113] = 32'h0;  // 32'h1de811e0;
    ram_cell[     114] = 32'h0;  // 32'hc524f2c6;
    ram_cell[     115] = 32'h0;  // 32'h03f20edc;
    ram_cell[     116] = 32'h0;  // 32'h2f05ac7f;
    ram_cell[     117] = 32'h0;  // 32'h71adec90;
    ram_cell[     118] = 32'h0;  // 32'ha3d54f7e;
    ram_cell[     119] = 32'h0;  // 32'hded935ad;
    ram_cell[     120] = 32'h0;  // 32'h9b4fee81;
    ram_cell[     121] = 32'h0;  // 32'hd49d6b0b;
    ram_cell[     122] = 32'h0;  // 32'hf286a429;
    ram_cell[     123] = 32'h0;  // 32'h997e2e44;
    ram_cell[     124] = 32'h0;  // 32'h32345b74;
    ram_cell[     125] = 32'h0;  // 32'hff3892b5;
    ram_cell[     126] = 32'h0;  // 32'h421d284f;
    ram_cell[     127] = 32'h0;  // 32'hfbaa48a7;
    ram_cell[     128] = 32'h0;  // 32'h9eed6bf1;
    ram_cell[     129] = 32'h0;  // 32'hfca3fd26;
    ram_cell[     130] = 32'h0;  // 32'h197ff06d;
    ram_cell[     131] = 32'h0;  // 32'h5ab06ebc;
    ram_cell[     132] = 32'h0;  // 32'h956c4efb;
    ram_cell[     133] = 32'h0;  // 32'hd60a1d6c;
    ram_cell[     134] = 32'h0;  // 32'he64caf81;
    ram_cell[     135] = 32'h0;  // 32'hca840497;
    ram_cell[     136] = 32'h0;  // 32'h1172fb5a;
    ram_cell[     137] = 32'h0;  // 32'hc976ab35;
    ram_cell[     138] = 32'h0;  // 32'h97b7d491;
    ram_cell[     139] = 32'h0;  // 32'he1e97ea4;
    ram_cell[     140] = 32'h0;  // 32'h579a607b;
    ram_cell[     141] = 32'h0;  // 32'hd055d0f4;
    ram_cell[     142] = 32'h0;  // 32'hdc2344f1;
    ram_cell[     143] = 32'h0;  // 32'h47ae4c2f;
    ram_cell[     144] = 32'h0;  // 32'h9a982947;
    ram_cell[     145] = 32'h0;  // 32'h1f6e210f;
    ram_cell[     146] = 32'h0;  // 32'hac6f68b7;
    ram_cell[     147] = 32'h0;  // 32'h7d0ba9be;
    ram_cell[     148] = 32'h0;  // 32'hc0b74b74;
    ram_cell[     149] = 32'h0;  // 32'h053b1bf4;
    ram_cell[     150] = 32'h0;  // 32'hce23fb73;
    ram_cell[     151] = 32'h0;  // 32'h83596f0f;
    ram_cell[     152] = 32'h0;  // 32'ha7ea217e;
    ram_cell[     153] = 32'h0;  // 32'h771c080b;
    ram_cell[     154] = 32'h0;  // 32'h3c1147cc;
    ram_cell[     155] = 32'h0;  // 32'hbf1f8406;
    ram_cell[     156] = 32'h0;  // 32'hf8a22518;
    ram_cell[     157] = 32'h0;  // 32'hf5319ad0;
    ram_cell[     158] = 32'h0;  // 32'hbf9f6217;
    ram_cell[     159] = 32'h0;  // 32'haf1e6f66;
    ram_cell[     160] = 32'h0;  // 32'h3c786e6d;
    ram_cell[     161] = 32'h0;  // 32'h7dec66bf;
    ram_cell[     162] = 32'h0;  // 32'h8336b9d7;
    ram_cell[     163] = 32'h0;  // 32'hde83b9f9;
    ram_cell[     164] = 32'h0;  // 32'h94dbcfb2;
    ram_cell[     165] = 32'h0;  // 32'h335283ec;
    ram_cell[     166] = 32'h0;  // 32'h2e349a82;
    ram_cell[     167] = 32'h0;  // 32'h360e2be1;
    ram_cell[     168] = 32'h0;  // 32'h0e8dc748;
    ram_cell[     169] = 32'h0;  // 32'h89e4a02e;
    ram_cell[     170] = 32'h0;  // 32'h0b3d2411;
    ram_cell[     171] = 32'h0;  // 32'hf9a67e65;
    ram_cell[     172] = 32'h0;  // 32'h0f72c681;
    ram_cell[     173] = 32'h0;  // 32'hf8800778;
    ram_cell[     174] = 32'h0;  // 32'h7c6b8916;
    ram_cell[     175] = 32'h0;  // 32'h31588076;
    ram_cell[     176] = 32'h0;  // 32'h30fd5c59;
    ram_cell[     177] = 32'h0;  // 32'h9cee5410;
    ram_cell[     178] = 32'h0;  // 32'h74494002;
    ram_cell[     179] = 32'h0;  // 32'h89ea9e77;
    ram_cell[     180] = 32'h0;  // 32'h97219ffc;
    ram_cell[     181] = 32'h0;  // 32'h37f44235;
    ram_cell[     182] = 32'h0;  // 32'h3e9012ed;
    ram_cell[     183] = 32'h0;  // 32'h52054a82;
    ram_cell[     184] = 32'h0;  // 32'ha1cb40c6;
    ram_cell[     185] = 32'h0;  // 32'h41e60b3f;
    ram_cell[     186] = 32'h0;  // 32'hf0167d38;
    ram_cell[     187] = 32'h0;  // 32'h642b08f1;
    ram_cell[     188] = 32'h0;  // 32'h55c36c16;
    ram_cell[     189] = 32'h0;  // 32'h63a8eefe;
    ram_cell[     190] = 32'h0;  // 32'h06a79a97;
    ram_cell[     191] = 32'h0;  // 32'h829a6979;
    ram_cell[     192] = 32'h0;  // 32'h958108f2;
    ram_cell[     193] = 32'h0;  // 32'h31d1ab7a;
    ram_cell[     194] = 32'h0;  // 32'h89695fcf;
    ram_cell[     195] = 32'h0;  // 32'h1a716cda;
    ram_cell[     196] = 32'h0;  // 32'hc09de17a;
    ram_cell[     197] = 32'h0;  // 32'h5b1d3524;
    ram_cell[     198] = 32'h0;  // 32'hd18cfc0c;
    ram_cell[     199] = 32'h0;  // 32'hf4350564;
    ram_cell[     200] = 32'h0;  // 32'h6a00d2e4;
    ram_cell[     201] = 32'h0;  // 32'h47a802bb;
    ram_cell[     202] = 32'h0;  // 32'hcd794b53;
    ram_cell[     203] = 32'h0;  // 32'h799e8658;
    ram_cell[     204] = 32'h0;  // 32'had4656bf;
    ram_cell[     205] = 32'h0;  // 32'hb027fabc;
    ram_cell[     206] = 32'h0;  // 32'hce79aa9b;
    ram_cell[     207] = 32'h0;  // 32'h758948fc;
    ram_cell[     208] = 32'h0;  // 32'h2678262c;
    ram_cell[     209] = 32'h0;  // 32'h13bca7a0;
    ram_cell[     210] = 32'h0;  // 32'h5ac02f61;
    ram_cell[     211] = 32'h0;  // 32'h7f81fffb;
    ram_cell[     212] = 32'h0;  // 32'he7c3f07d;
    ram_cell[     213] = 32'h0;  // 32'he03cf28a;
    ram_cell[     214] = 32'h0;  // 32'h9b1968fc;
    ram_cell[     215] = 32'h0;  // 32'h79ee27ea;
    ram_cell[     216] = 32'h0;  // 32'ha6850ab3;
    ram_cell[     217] = 32'h0;  // 32'h89b8fc7a;
    ram_cell[     218] = 32'h0;  // 32'h6a5c1199;
    ram_cell[     219] = 32'h0;  // 32'h89c9c143;
    ram_cell[     220] = 32'h0;  // 32'h831cd878;
    ram_cell[     221] = 32'h0;  // 32'hb17b7deb;
    ram_cell[     222] = 32'h0;  // 32'h6b761676;
    ram_cell[     223] = 32'h0;  // 32'h01ee4f4b;
    ram_cell[     224] = 32'h0;  // 32'h53c1a7ed;
    ram_cell[     225] = 32'h0;  // 32'heb584f94;
    ram_cell[     226] = 32'h0;  // 32'hc7441873;
    ram_cell[     227] = 32'h0;  // 32'h1f627fe1;
    ram_cell[     228] = 32'h0;  // 32'h8e4b66d7;
    ram_cell[     229] = 32'h0;  // 32'h81ff60b9;
    ram_cell[     230] = 32'h0;  // 32'hd816051a;
    ram_cell[     231] = 32'h0;  // 32'hdd71af83;
    ram_cell[     232] = 32'h0;  // 32'hb879040e;
    ram_cell[     233] = 32'h0;  // 32'ha81179f5;
    ram_cell[     234] = 32'h0;  // 32'h1bb91d31;
    ram_cell[     235] = 32'h0;  // 32'hc9150244;
    ram_cell[     236] = 32'h0;  // 32'hf73c8757;
    ram_cell[     237] = 32'h0;  // 32'h90febc77;
    ram_cell[     238] = 32'h0;  // 32'ha4b97d01;
    ram_cell[     239] = 32'h0;  // 32'h1e1f0689;
    ram_cell[     240] = 32'h0;  // 32'heb37fb2b;
    ram_cell[     241] = 32'h0;  // 32'h783f9fe5;
    ram_cell[     242] = 32'h0;  // 32'h380f6401;
    ram_cell[     243] = 32'h0;  // 32'h1fb73a27;
    ram_cell[     244] = 32'h0;  // 32'h9a4a3845;
    ram_cell[     245] = 32'h0;  // 32'hab911604;
    ram_cell[     246] = 32'h0;  // 32'hdc353444;
    ram_cell[     247] = 32'h0;  // 32'hf461a96e;
    ram_cell[     248] = 32'h0;  // 32'h36474898;
    ram_cell[     249] = 32'h0;  // 32'h11eaab79;
    ram_cell[     250] = 32'h0;  // 32'h7b886261;
    ram_cell[     251] = 32'h0;  // 32'h30806ac7;
    ram_cell[     252] = 32'h0;  // 32'h7796a478;
    ram_cell[     253] = 32'h0;  // 32'he99bef5a;
    ram_cell[     254] = 32'h0;  // 32'h7e6fe510;
    ram_cell[     255] = 32'h0;  // 32'h662d418c;
    // src matrix A
    ram_cell[     256] = 32'h6170d581;
    ram_cell[     257] = 32'h3b935766;
    ram_cell[     258] = 32'h6bb6d245;
    ram_cell[     259] = 32'h8808a48e;
    ram_cell[     260] = 32'h37c1a9e0;
    ram_cell[     261] = 32'haa7ae776;
    ram_cell[     262] = 32'hb7ff5685;
    ram_cell[     263] = 32'he3174a69;
    ram_cell[     264] = 32'hfd2756b0;
    ram_cell[     265] = 32'hc8d9cc3d;
    ram_cell[     266] = 32'hef085bb6;
    ram_cell[     267] = 32'hdb39a9d5;
    ram_cell[     268] = 32'h523a40ff;
    ram_cell[     269] = 32'h7c6c6802;
    ram_cell[     270] = 32'hf39c87d9;
    ram_cell[     271] = 32'h51cbf7a5;
    ram_cell[     272] = 32'h6b4fcf52;
    ram_cell[     273] = 32'h4d2fa379;
    ram_cell[     274] = 32'h18e43b92;
    ram_cell[     275] = 32'h9beac867;
    ram_cell[     276] = 32'h33e202a3;
    ram_cell[     277] = 32'h0e06b208;
    ram_cell[     278] = 32'h36a1c04c;
    ram_cell[     279] = 32'he66da79a;
    ram_cell[     280] = 32'h642f0930;
    ram_cell[     281] = 32'h242d5c28;
    ram_cell[     282] = 32'hc9eb0864;
    ram_cell[     283] = 32'h4900e337;
    ram_cell[     284] = 32'hcabd403d;
    ram_cell[     285] = 32'h52088362;
    ram_cell[     286] = 32'h0b88bfa7;
    ram_cell[     287] = 32'h04c0f833;
    ram_cell[     288] = 32'hdcbc239b;
    ram_cell[     289] = 32'h04170112;
    ram_cell[     290] = 32'h209291a8;
    ram_cell[     291] = 32'hccaa3fa0;
    ram_cell[     292] = 32'h8d177aa7;
    ram_cell[     293] = 32'hd97c1fc2;
    ram_cell[     294] = 32'hc8b1dfbf;
    ram_cell[     295] = 32'h2091d0f6;
    ram_cell[     296] = 32'h13e7fbe6;
    ram_cell[     297] = 32'hf8ee11cf;
    ram_cell[     298] = 32'ha6c801f1;
    ram_cell[     299] = 32'hd1db9121;
    ram_cell[     300] = 32'h1bfcfb92;
    ram_cell[     301] = 32'h182adf8e;
    ram_cell[     302] = 32'h366984ae;
    ram_cell[     303] = 32'hd4284a6a;
    ram_cell[     304] = 32'hce4b4539;
    ram_cell[     305] = 32'h6c8fba8c;
    ram_cell[     306] = 32'h22c5bf20;
    ram_cell[     307] = 32'h9b87682e;
    ram_cell[     308] = 32'h97db7948;
    ram_cell[     309] = 32'h9cd0eefa;
    ram_cell[     310] = 32'h7d343d4b;
    ram_cell[     311] = 32'hc5052548;
    ram_cell[     312] = 32'h274a3bc2;
    ram_cell[     313] = 32'h0eb5429f;
    ram_cell[     314] = 32'heb5980ea;
    ram_cell[     315] = 32'h7004aa97;
    ram_cell[     316] = 32'hacdd3cfe;
    ram_cell[     317] = 32'h526d4040;
    ram_cell[     318] = 32'hc3f8fc34;
    ram_cell[     319] = 32'h3407e9ab;
    ram_cell[     320] = 32'h490376cd;
    ram_cell[     321] = 32'h2ed13fbb;
    ram_cell[     322] = 32'hc8e684d8;
    ram_cell[     323] = 32'he5e9d30c;
    ram_cell[     324] = 32'hccaa4d56;
    ram_cell[     325] = 32'hd589ef13;
    ram_cell[     326] = 32'h507e1e7c;
    ram_cell[     327] = 32'h2b4a2699;
    ram_cell[     328] = 32'h289b2568;
    ram_cell[     329] = 32'h8e89cfac;
    ram_cell[     330] = 32'h902bda30;
    ram_cell[     331] = 32'h3b5d0c3b;
    ram_cell[     332] = 32'h1b1e549b;
    ram_cell[     333] = 32'hc22fe87a;
    ram_cell[     334] = 32'hf6fd2c2b;
    ram_cell[     335] = 32'had09715b;
    ram_cell[     336] = 32'hf3710f94;
    ram_cell[     337] = 32'hddfd4420;
    ram_cell[     338] = 32'hd7ffd29b;
    ram_cell[     339] = 32'hb83c49e9;
    ram_cell[     340] = 32'h324b6e47;
    ram_cell[     341] = 32'h0a950a40;
    ram_cell[     342] = 32'h2412f5ec;
    ram_cell[     343] = 32'he840b37a;
    ram_cell[     344] = 32'h10133c63;
    ram_cell[     345] = 32'h3e2c5fba;
    ram_cell[     346] = 32'hb0c0c0e1;
    ram_cell[     347] = 32'h8dff54f5;
    ram_cell[     348] = 32'h96788167;
    ram_cell[     349] = 32'hf1bff0f4;
    ram_cell[     350] = 32'h6f05d8eb;
    ram_cell[     351] = 32'h56e266d6;
    ram_cell[     352] = 32'h42f1d140;
    ram_cell[     353] = 32'h1a00db35;
    ram_cell[     354] = 32'h5b085907;
    ram_cell[     355] = 32'h0a6541ad;
    ram_cell[     356] = 32'h12fa1844;
    ram_cell[     357] = 32'h8d3f804a;
    ram_cell[     358] = 32'h361d9e2f;
    ram_cell[     359] = 32'h4e200aa8;
    ram_cell[     360] = 32'hab2b3e38;
    ram_cell[     361] = 32'h391a1152;
    ram_cell[     362] = 32'hf2667916;
    ram_cell[     363] = 32'h1906e817;
    ram_cell[     364] = 32'hab06e590;
    ram_cell[     365] = 32'h0bd56fd8;
    ram_cell[     366] = 32'h569d7f26;
    ram_cell[     367] = 32'h78adff87;
    ram_cell[     368] = 32'h6cffba6a;
    ram_cell[     369] = 32'hda6064e0;
    ram_cell[     370] = 32'h5aa8be79;
    ram_cell[     371] = 32'h5dc0e2b8;
    ram_cell[     372] = 32'h9483e9c5;
    ram_cell[     373] = 32'h40854240;
    ram_cell[     374] = 32'h0dbba311;
    ram_cell[     375] = 32'hdeab299f;
    ram_cell[     376] = 32'h608c4edc;
    ram_cell[     377] = 32'hea53f1b2;
    ram_cell[     378] = 32'h1787c573;
    ram_cell[     379] = 32'hea969c51;
    ram_cell[     380] = 32'h43b91742;
    ram_cell[     381] = 32'hb51258f1;
    ram_cell[     382] = 32'h4ca0edeb;
    ram_cell[     383] = 32'h58f9233d;
    ram_cell[     384] = 32'h81fc63a8;
    ram_cell[     385] = 32'hce16a6a3;
    ram_cell[     386] = 32'h66a79caf;
    ram_cell[     387] = 32'hba372498;
    ram_cell[     388] = 32'hf942812e;
    ram_cell[     389] = 32'h8c431a09;
    ram_cell[     390] = 32'hcae01a51;
    ram_cell[     391] = 32'hffe1a436;
    ram_cell[     392] = 32'h88bab75a;
    ram_cell[     393] = 32'h6338dafa;
    ram_cell[     394] = 32'h77af5af9;
    ram_cell[     395] = 32'h14de4a5b;
    ram_cell[     396] = 32'h428e6920;
    ram_cell[     397] = 32'h740869db;
    ram_cell[     398] = 32'hca65ec9d;
    ram_cell[     399] = 32'hdf18002a;
    ram_cell[     400] = 32'h05e5f659;
    ram_cell[     401] = 32'h64e114db;
    ram_cell[     402] = 32'h0ff5ab1c;
    ram_cell[     403] = 32'h2f54a4fc;
    ram_cell[     404] = 32'h27438d00;
    ram_cell[     405] = 32'hfb49d7bf;
    ram_cell[     406] = 32'h6f8bedcc;
    ram_cell[     407] = 32'h7c33f629;
    ram_cell[     408] = 32'hc9f0aad8;
    ram_cell[     409] = 32'h5cefe3d9;
    ram_cell[     410] = 32'hf798bdb2;
    ram_cell[     411] = 32'h11bc7dc6;
    ram_cell[     412] = 32'h1520cd52;
    ram_cell[     413] = 32'hf032c5f5;
    ram_cell[     414] = 32'hcceb230b;
    ram_cell[     415] = 32'ha29427fc;
    ram_cell[     416] = 32'hdeeeede7;
    ram_cell[     417] = 32'hd7a5de9e;
    ram_cell[     418] = 32'h7c9d9a92;
    ram_cell[     419] = 32'h099504f7;
    ram_cell[     420] = 32'hc733463e;
    ram_cell[     421] = 32'h78842a2f;
    ram_cell[     422] = 32'h3ef0accd;
    ram_cell[     423] = 32'h8850a0b5;
    ram_cell[     424] = 32'h23528d69;
    ram_cell[     425] = 32'h41c7eb9e;
    ram_cell[     426] = 32'he096918b;
    ram_cell[     427] = 32'h99111f03;
    ram_cell[     428] = 32'he6cbc849;
    ram_cell[     429] = 32'h7b99875b;
    ram_cell[     430] = 32'h11e0ed78;
    ram_cell[     431] = 32'ha693cc91;
    ram_cell[     432] = 32'ha1aadb76;
    ram_cell[     433] = 32'hb472a594;
    ram_cell[     434] = 32'hcfb78ad8;
    ram_cell[     435] = 32'hd72b058f;
    ram_cell[     436] = 32'hb06fa89f;
    ram_cell[     437] = 32'h6fe1b31f;
    ram_cell[     438] = 32'hdb90b49e;
    ram_cell[     439] = 32'h805509c2;
    ram_cell[     440] = 32'h8ca9286d;
    ram_cell[     441] = 32'hc96b0fa0;
    ram_cell[     442] = 32'he4f1f74c;
    ram_cell[     443] = 32'h464c9382;
    ram_cell[     444] = 32'h9bc41be9;
    ram_cell[     445] = 32'h23f8c9c6;
    ram_cell[     446] = 32'hf64756ec;
    ram_cell[     447] = 32'h4e5d58c2;
    ram_cell[     448] = 32'h53bbfbb1;
    ram_cell[     449] = 32'hbdd0ccff;
    ram_cell[     450] = 32'hb385ceec;
    ram_cell[     451] = 32'h4dc70063;
    ram_cell[     452] = 32'he80851c3;
    ram_cell[     453] = 32'he0d00ac1;
    ram_cell[     454] = 32'h4ed1736c;
    ram_cell[     455] = 32'h7738ec63;
    ram_cell[     456] = 32'hade58067;
    ram_cell[     457] = 32'h114b47d3;
    ram_cell[     458] = 32'hf2ff82fa;
    ram_cell[     459] = 32'h021c2246;
    ram_cell[     460] = 32'hc1fcf0bf;
    ram_cell[     461] = 32'h20e0b740;
    ram_cell[     462] = 32'h8f65bf09;
    ram_cell[     463] = 32'ha6e2b590;
    ram_cell[     464] = 32'h0387d72a;
    ram_cell[     465] = 32'h2809cb12;
    ram_cell[     466] = 32'hed8f3ea4;
    ram_cell[     467] = 32'hdf582ae8;
    ram_cell[     468] = 32'hb94b2d45;
    ram_cell[     469] = 32'h9c02577f;
    ram_cell[     470] = 32'hb6fab27f;
    ram_cell[     471] = 32'h31644696;
    ram_cell[     472] = 32'hb58e2c2f;
    ram_cell[     473] = 32'h5c951332;
    ram_cell[     474] = 32'h44fb2156;
    ram_cell[     475] = 32'h813eb46b;
    ram_cell[     476] = 32'hf3f4cac1;
    ram_cell[     477] = 32'h97637fe8;
    ram_cell[     478] = 32'h3d6f5cf1;
    ram_cell[     479] = 32'h7c76e352;
    ram_cell[     480] = 32'h4ea641eb;
    ram_cell[     481] = 32'h480a5ee2;
    ram_cell[     482] = 32'h7add1e09;
    ram_cell[     483] = 32'h2e49a57c;
    ram_cell[     484] = 32'h9915a25b;
    ram_cell[     485] = 32'he30b1de6;
    ram_cell[     486] = 32'h8605c1e2;
    ram_cell[     487] = 32'hb8363b8e;
    ram_cell[     488] = 32'ha6d82620;
    ram_cell[     489] = 32'h2b4c3f54;
    ram_cell[     490] = 32'h534c76fe;
    ram_cell[     491] = 32'ha8bca954;
    ram_cell[     492] = 32'he5c7d882;
    ram_cell[     493] = 32'h97bceb5a;
    ram_cell[     494] = 32'hb20fcdf4;
    ram_cell[     495] = 32'h897cdd20;
    ram_cell[     496] = 32'h6ed4c596;
    ram_cell[     497] = 32'h1187cba3;
    ram_cell[     498] = 32'h6b7adc52;
    ram_cell[     499] = 32'hb011f7b8;
    ram_cell[     500] = 32'h05f3207b;
    ram_cell[     501] = 32'h898a57c7;
    ram_cell[     502] = 32'ha04ad974;
    ram_cell[     503] = 32'hef19b7c1;
    ram_cell[     504] = 32'h646757fb;
    ram_cell[     505] = 32'haabf2638;
    ram_cell[     506] = 32'h04f3fe59;
    ram_cell[     507] = 32'h0ab17f5b;
    ram_cell[     508] = 32'h013cd39c;
    ram_cell[     509] = 32'hfdc91374;
    ram_cell[     510] = 32'h90139f80;
    ram_cell[     511] = 32'hd68a532d;
    // src matrix B
    ram_cell[     512] = 32'h1182d9c9;
    ram_cell[     513] = 32'hf3b5cef6;
    ram_cell[     514] = 32'hfa1af7c9;
    ram_cell[     515] = 32'hc171a9d5;
    ram_cell[     516] = 32'hb0f34779;
    ram_cell[     517] = 32'h66eac363;
    ram_cell[     518] = 32'h85cae939;
    ram_cell[     519] = 32'h632f1559;
    ram_cell[     520] = 32'h89220de3;
    ram_cell[     521] = 32'hdc6c3bef;
    ram_cell[     522] = 32'ha909c551;
    ram_cell[     523] = 32'h82009fe5;
    ram_cell[     524] = 32'h1de5b42e;
    ram_cell[     525] = 32'h769eacfd;
    ram_cell[     526] = 32'h35d4821f;
    ram_cell[     527] = 32'hdfc90079;
    ram_cell[     528] = 32'h134eaa9a;
    ram_cell[     529] = 32'h0817d80a;
    ram_cell[     530] = 32'haf70bc1c;
    ram_cell[     531] = 32'he226ba80;
    ram_cell[     532] = 32'h458cdd01;
    ram_cell[     533] = 32'hd37042e2;
    ram_cell[     534] = 32'hfa7a689d;
    ram_cell[     535] = 32'h48daace6;
    ram_cell[     536] = 32'h68de8f2f;
    ram_cell[     537] = 32'h4039ca30;
    ram_cell[     538] = 32'h30fda0c0;
    ram_cell[     539] = 32'hab956e0e;
    ram_cell[     540] = 32'hb15b8ac1;
    ram_cell[     541] = 32'h3a8824e7;
    ram_cell[     542] = 32'ha1a845a9;
    ram_cell[     543] = 32'h2ce763e7;
    ram_cell[     544] = 32'hf7c636fe;
    ram_cell[     545] = 32'h4a2bacf3;
    ram_cell[     546] = 32'h22da56f6;
    ram_cell[     547] = 32'hff83299c;
    ram_cell[     548] = 32'h58519bff;
    ram_cell[     549] = 32'h09e53a7a;
    ram_cell[     550] = 32'h988f897f;
    ram_cell[     551] = 32'h6acbb1f8;
    ram_cell[     552] = 32'hda084552;
    ram_cell[     553] = 32'h501024be;
    ram_cell[     554] = 32'h65d28b87;
    ram_cell[     555] = 32'h2263f6f3;
    ram_cell[     556] = 32'h019982d0;
    ram_cell[     557] = 32'h13dec7a3;
    ram_cell[     558] = 32'h297534f5;
    ram_cell[     559] = 32'h410acf12;
    ram_cell[     560] = 32'h0be03b6b;
    ram_cell[     561] = 32'h8d9bde87;
    ram_cell[     562] = 32'h538a721b;
    ram_cell[     563] = 32'h91648b31;
    ram_cell[     564] = 32'h87a34d07;
    ram_cell[     565] = 32'h59be7edc;
    ram_cell[     566] = 32'h977dc66d;
    ram_cell[     567] = 32'hd72c3d73;
    ram_cell[     568] = 32'h89e24d71;
    ram_cell[     569] = 32'h880caff8;
    ram_cell[     570] = 32'h968366b6;
    ram_cell[     571] = 32'hb23bb8d3;
    ram_cell[     572] = 32'hab3c3752;
    ram_cell[     573] = 32'h8245f066;
    ram_cell[     574] = 32'h399f9957;
    ram_cell[     575] = 32'h6a1e8c60;
    ram_cell[     576] = 32'hb1df0b4e;
    ram_cell[     577] = 32'hc523fedb;
    ram_cell[     578] = 32'h850a8600;
    ram_cell[     579] = 32'hc90c6f48;
    ram_cell[     580] = 32'h3513c231;
    ram_cell[     581] = 32'he32f09b0;
    ram_cell[     582] = 32'h32bb92f2;
    ram_cell[     583] = 32'h6f6412ee;
    ram_cell[     584] = 32'hf1edafb3;
    ram_cell[     585] = 32'hfe8bf804;
    ram_cell[     586] = 32'h5706b879;
    ram_cell[     587] = 32'heb187b42;
    ram_cell[     588] = 32'h0b4ad82b;
    ram_cell[     589] = 32'hfddb67e5;
    ram_cell[     590] = 32'h19ae574b;
    ram_cell[     591] = 32'hf43c31b4;
    ram_cell[     592] = 32'h34bfcb99;
    ram_cell[     593] = 32'h818f6824;
    ram_cell[     594] = 32'h9d269ac9;
    ram_cell[     595] = 32'hd6bba0ad;
    ram_cell[     596] = 32'hbf57c153;
    ram_cell[     597] = 32'hd40708fb;
    ram_cell[     598] = 32'h75cc5580;
    ram_cell[     599] = 32'hea5bc862;
    ram_cell[     600] = 32'h8e985495;
    ram_cell[     601] = 32'h0ce4d7f8;
    ram_cell[     602] = 32'h22e21d99;
    ram_cell[     603] = 32'h4982f11b;
    ram_cell[     604] = 32'hf3b54543;
    ram_cell[     605] = 32'h4b533b0a;
    ram_cell[     606] = 32'h1655c69d;
    ram_cell[     607] = 32'h43e4a5a7;
    ram_cell[     608] = 32'h1e0d0ea2;
    ram_cell[     609] = 32'h860e6d61;
    ram_cell[     610] = 32'h58f54f19;
    ram_cell[     611] = 32'h88d786ea;
    ram_cell[     612] = 32'h426d9938;
    ram_cell[     613] = 32'hbf7755ed;
    ram_cell[     614] = 32'hb43216b8;
    ram_cell[     615] = 32'hc64f5141;
    ram_cell[     616] = 32'h0aa14608;
    ram_cell[     617] = 32'h11123cfa;
    ram_cell[     618] = 32'hede0f70e;
    ram_cell[     619] = 32'hfc0e28c5;
    ram_cell[     620] = 32'h20bac925;
    ram_cell[     621] = 32'ha7f30bc4;
    ram_cell[     622] = 32'hb829b0d7;
    ram_cell[     623] = 32'h4e60023c;
    ram_cell[     624] = 32'h0ae5f060;
    ram_cell[     625] = 32'hcf90898e;
    ram_cell[     626] = 32'h640978da;
    ram_cell[     627] = 32'hc8ade098;
    ram_cell[     628] = 32'h8240f8e9;
    ram_cell[     629] = 32'h805bb9de;
    ram_cell[     630] = 32'h68cce09a;
    ram_cell[     631] = 32'he58414d1;
    ram_cell[     632] = 32'h6784c54d;
    ram_cell[     633] = 32'h339f5ecf;
    ram_cell[     634] = 32'h6cbecaea;
    ram_cell[     635] = 32'h2660ee25;
    ram_cell[     636] = 32'h98a59eda;
    ram_cell[     637] = 32'h119a2801;
    ram_cell[     638] = 32'h1b4e982a;
    ram_cell[     639] = 32'hd974ee34;
    ram_cell[     640] = 32'h1710994e;
    ram_cell[     641] = 32'h39f59da4;
    ram_cell[     642] = 32'hbf474384;
    ram_cell[     643] = 32'heac969c7;
    ram_cell[     644] = 32'h9ec37843;
    ram_cell[     645] = 32'hf9fc64b0;
    ram_cell[     646] = 32'h06c148d3;
    ram_cell[     647] = 32'h29a3f2ae;
    ram_cell[     648] = 32'ha667a8bc;
    ram_cell[     649] = 32'hf52f4920;
    ram_cell[     650] = 32'h54140434;
    ram_cell[     651] = 32'h7a95f2ea;
    ram_cell[     652] = 32'he119b0b0;
    ram_cell[     653] = 32'h92167d0c;
    ram_cell[     654] = 32'h74ae9bc3;
    ram_cell[     655] = 32'hd8aec3c8;
    ram_cell[     656] = 32'had3cad01;
    ram_cell[     657] = 32'h83ed608c;
    ram_cell[     658] = 32'h72c75c58;
    ram_cell[     659] = 32'h0898459b;
    ram_cell[     660] = 32'h5aec9de0;
    ram_cell[     661] = 32'hf711bd86;
    ram_cell[     662] = 32'he372a9ee;
    ram_cell[     663] = 32'h5469bf4b;
    ram_cell[     664] = 32'he8cef907;
    ram_cell[     665] = 32'hfa018adb;
    ram_cell[     666] = 32'hbc51ab6a;
    ram_cell[     667] = 32'hd2f54ee9;
    ram_cell[     668] = 32'h2443ffa5;
    ram_cell[     669] = 32'hc2dd62bc;
    ram_cell[     670] = 32'hae57ddd6;
    ram_cell[     671] = 32'h020b2734;
    ram_cell[     672] = 32'h3b83bb85;
    ram_cell[     673] = 32'h80e3c2eb;
    ram_cell[     674] = 32'hd416ed05;
    ram_cell[     675] = 32'h5a794094;
    ram_cell[     676] = 32'haff6dc31;
    ram_cell[     677] = 32'hee7faef2;
    ram_cell[     678] = 32'haf93a44d;
    ram_cell[     679] = 32'ha73f995b;
    ram_cell[     680] = 32'hc581411b;
    ram_cell[     681] = 32'h845302b3;
    ram_cell[     682] = 32'h6c913a3c;
    ram_cell[     683] = 32'h70e13f17;
    ram_cell[     684] = 32'h5e612ec9;
    ram_cell[     685] = 32'ha6c4b54f;
    ram_cell[     686] = 32'h56bc0f12;
    ram_cell[     687] = 32'h78965b6b;
    ram_cell[     688] = 32'h35361411;
    ram_cell[     689] = 32'ha27a4a66;
    ram_cell[     690] = 32'h5940d345;
    ram_cell[     691] = 32'h6cc47b0e;
    ram_cell[     692] = 32'h5d7e6d21;
    ram_cell[     693] = 32'h76c26c62;
    ram_cell[     694] = 32'hd7c5195f;
    ram_cell[     695] = 32'hae0973db;
    ram_cell[     696] = 32'hf6a32eda;
    ram_cell[     697] = 32'hb0e7ab72;
    ram_cell[     698] = 32'h1f5723d5;
    ram_cell[     699] = 32'hf2de532a;
    ram_cell[     700] = 32'hf08de3ba;
    ram_cell[     701] = 32'h98d34254;
    ram_cell[     702] = 32'h6cbdef09;
    ram_cell[     703] = 32'h760b6c2b;
    ram_cell[     704] = 32'h9cfe2e3d;
    ram_cell[     705] = 32'h502f399c;
    ram_cell[     706] = 32'hc6db5420;
    ram_cell[     707] = 32'h07dac942;
    ram_cell[     708] = 32'h1ed48dda;
    ram_cell[     709] = 32'h72993f5c;
    ram_cell[     710] = 32'h62c774a1;
    ram_cell[     711] = 32'hec4fe1d9;
    ram_cell[     712] = 32'hf91e4893;
    ram_cell[     713] = 32'h137b2e7b;
    ram_cell[     714] = 32'h5a576a7a;
    ram_cell[     715] = 32'hca9b4697;
    ram_cell[     716] = 32'hd9ccd606;
    ram_cell[     717] = 32'h23bbf9a1;
    ram_cell[     718] = 32'hba369d69;
    ram_cell[     719] = 32'h477300a2;
    ram_cell[     720] = 32'h5ce02163;
    ram_cell[     721] = 32'h7acc9169;
    ram_cell[     722] = 32'h30c4d381;
    ram_cell[     723] = 32'h13aea518;
    ram_cell[     724] = 32'h7e897445;
    ram_cell[     725] = 32'hc957108a;
    ram_cell[     726] = 32'hb7179d7c;
    ram_cell[     727] = 32'ha06a611b;
    ram_cell[     728] = 32'hcf3c0f13;
    ram_cell[     729] = 32'h431b7ee3;
    ram_cell[     730] = 32'ha6a55204;
    ram_cell[     731] = 32'hc32ee114;
    ram_cell[     732] = 32'hf3ccfce8;
    ram_cell[     733] = 32'h2f700b5e;
    ram_cell[     734] = 32'hb023d660;
    ram_cell[     735] = 32'h125fb370;
    ram_cell[     736] = 32'hda3933d1;
    ram_cell[     737] = 32'h23220e2c;
    ram_cell[     738] = 32'h751b8898;
    ram_cell[     739] = 32'h1f1dab33;
    ram_cell[     740] = 32'h08baf117;
    ram_cell[     741] = 32'h975db85a;
    ram_cell[     742] = 32'haf047447;
    ram_cell[     743] = 32'h68cb37d3;
    ram_cell[     744] = 32'hb97e51b4;
    ram_cell[     745] = 32'h4c340765;
    ram_cell[     746] = 32'h1bc1cba4;
    ram_cell[     747] = 32'hb2dae800;
    ram_cell[     748] = 32'h7a178cc3;
    ram_cell[     749] = 32'h0b2f769f;
    ram_cell[     750] = 32'haff59dc2;
    ram_cell[     751] = 32'h6eebabbd;
    ram_cell[     752] = 32'hf92b7d6e;
    ram_cell[     753] = 32'h77d73e4d;
    ram_cell[     754] = 32'h1cfcf1ec;
    ram_cell[     755] = 32'ha62f97e1;
    ram_cell[     756] = 32'h27d209ec;
    ram_cell[     757] = 32'h3f2bc993;
    ram_cell[     758] = 32'h4ab3c1d4;
    ram_cell[     759] = 32'hd7025503;
    ram_cell[     760] = 32'h6874bc7f;
    ram_cell[     761] = 32'h8868a515;
    ram_cell[     762] = 32'h90d24d94;
    ram_cell[     763] = 32'h73aa6d12;
    ram_cell[     764] = 32'h07488ae8;
    ram_cell[     765] = 32'h81bb283e;
    ram_cell[     766] = 32'h27016d41;
    ram_cell[     767] = 32'hb0bc3290;
end

endmodule

