module bht(
    
);

endmodule