
module mem #(                   // 
    parameter  ADDR_LEN  = 11   // 
) (
    input  clk, rst,
    input  [ADDR_LEN-1:0] addr, // memory address
    output reg [31:0] rd_data,  // data read out
    input  wr_req,
    input  [31:0] wr_data       // data write in
);
localparam MEM_SIZE = 1<<ADDR_LEN;
reg [31:0] ram_cell [MEM_SIZE];

always @ (posedge clk or posedge rst)
    if(rst)
        rd_data <= 0;
    else
        rd_data <= ram_cell[addr];

always @ (posedge clk)
    if(wr_req) 
        ram_cell[addr] <= wr_data;

initial begin
    // dst matrix C
    ram_cell[       0] = 32'h0;  // 32'h378a25dd;
    ram_cell[       1] = 32'h0;  // 32'h1d52ed49;
    ram_cell[       2] = 32'h0;  // 32'h5ced846f;
    ram_cell[       3] = 32'h0;  // 32'h8b984e34;
    ram_cell[       4] = 32'h0;  // 32'h25ff5ceb;
    ram_cell[       5] = 32'h0;  // 32'h74da70e6;
    ram_cell[       6] = 32'h0;  // 32'h2521b465;
    ram_cell[       7] = 32'h0;  // 32'ha86787f0;
    ram_cell[       8] = 32'h0;  // 32'h47c70f83;
    ram_cell[       9] = 32'h0;  // 32'h730bfdb0;
    ram_cell[      10] = 32'h0;  // 32'h739e2839;
    ram_cell[      11] = 32'h0;  // 32'h24b8097f;
    ram_cell[      12] = 32'h0;  // 32'hae60d853;
    ram_cell[      13] = 32'h0;  // 32'h3e808252;
    ram_cell[      14] = 32'h0;  // 32'h211ea692;
    ram_cell[      15] = 32'h0;  // 32'hbd75bc4f;
    ram_cell[      16] = 32'h0;  // 32'h5e1dba0f;
    ram_cell[      17] = 32'h0;  // 32'hbda85daa;
    ram_cell[      18] = 32'h0;  // 32'hecb1bb85;
    ram_cell[      19] = 32'h0;  // 32'h3836fceb;
    ram_cell[      20] = 32'h0;  // 32'h58961ac6;
    ram_cell[      21] = 32'h0;  // 32'h75fb0a81;
    ram_cell[      22] = 32'h0;  // 32'hbe684008;
    ram_cell[      23] = 32'h0;  // 32'h5a903410;
    ram_cell[      24] = 32'h0;  // 32'hcc79d73a;
    ram_cell[      25] = 32'h0;  // 32'h8e75a337;
    ram_cell[      26] = 32'h0;  // 32'h80d4e2bf;
    ram_cell[      27] = 32'h0;  // 32'h40a88e94;
    ram_cell[      28] = 32'h0;  // 32'he0919ff9;
    ram_cell[      29] = 32'h0;  // 32'h94b27df9;
    ram_cell[      30] = 32'h0;  // 32'h257b4eb1;
    ram_cell[      31] = 32'h0;  // 32'ha975742f;
    ram_cell[      32] = 32'h0;  // 32'h1f5a89cd;
    ram_cell[      33] = 32'h0;  // 32'h0107701a;
    ram_cell[      34] = 32'h0;  // 32'h29579d50;
    ram_cell[      35] = 32'h0;  // 32'hb31d4e9e;
    ram_cell[      36] = 32'h0;  // 32'h25c23fc4;
    ram_cell[      37] = 32'h0;  // 32'h127d144b;
    ram_cell[      38] = 32'h0;  // 32'h5d70dc85;
    ram_cell[      39] = 32'h0;  // 32'h1215bcc9;
    ram_cell[      40] = 32'h0;  // 32'h67609af6;
    ram_cell[      41] = 32'h0;  // 32'h27e8d21f;
    ram_cell[      42] = 32'h0;  // 32'h79470eb8;
    ram_cell[      43] = 32'h0;  // 32'hb999e6d8;
    ram_cell[      44] = 32'h0;  // 32'h07ea4420;
    ram_cell[      45] = 32'h0;  // 32'ha486f445;
    ram_cell[      46] = 32'h0;  // 32'h8088ea1a;
    ram_cell[      47] = 32'h0;  // 32'h58273448;
    ram_cell[      48] = 32'h0;  // 32'hd6421441;
    ram_cell[      49] = 32'h0;  // 32'ha0e0a6a4;
    ram_cell[      50] = 32'h0;  // 32'h5d24e976;
    ram_cell[      51] = 32'h0;  // 32'h9c95b96d;
    ram_cell[      52] = 32'h0;  // 32'h3436cd1f;
    ram_cell[      53] = 32'h0;  // 32'h46c30e8b;
    ram_cell[      54] = 32'h0;  // 32'hb9883894;
    ram_cell[      55] = 32'h0;  // 32'h79016e48;
    ram_cell[      56] = 32'h0;  // 32'ha93f23e7;
    ram_cell[      57] = 32'h0;  // 32'he898577f;
    ram_cell[      58] = 32'h0;  // 32'h3daa3807;
    ram_cell[      59] = 32'h0;  // 32'hbce9c43b;
    ram_cell[      60] = 32'h0;  // 32'h56d726e4;
    ram_cell[      61] = 32'h0;  // 32'h73cfddc1;
    ram_cell[      62] = 32'h0;  // 32'h9138d9a5;
    ram_cell[      63] = 32'h0;  // 32'h9548bf9a;
    ram_cell[      64] = 32'h0;  // 32'h7a6a37f5;
    ram_cell[      65] = 32'h0;  // 32'ha089f344;
    ram_cell[      66] = 32'h0;  // 32'he98a5237;
    ram_cell[      67] = 32'h0;  // 32'hc760be80;
    ram_cell[      68] = 32'h0;  // 32'h24dee1d7;
    ram_cell[      69] = 32'h0;  // 32'h5279aec9;
    ram_cell[      70] = 32'h0;  // 32'hd463e7f7;
    ram_cell[      71] = 32'h0;  // 32'hea81d738;
    ram_cell[      72] = 32'h0;  // 32'h9bc10fbb;
    ram_cell[      73] = 32'h0;  // 32'h0b4c4096;
    ram_cell[      74] = 32'h0;  // 32'h112944b6;
    ram_cell[      75] = 32'h0;  // 32'h523e91e1;
    ram_cell[      76] = 32'h0;  // 32'h5c88872e;
    ram_cell[      77] = 32'h0;  // 32'h75feffa8;
    ram_cell[      78] = 32'h0;  // 32'h297363cf;
    ram_cell[      79] = 32'h0;  // 32'ha94d2a66;
    ram_cell[      80] = 32'h0;  // 32'h4e709bc9;
    ram_cell[      81] = 32'h0;  // 32'h13f0fd01;
    ram_cell[      82] = 32'h0;  // 32'h0e177e42;
    ram_cell[      83] = 32'h0;  // 32'h41f0be88;
    ram_cell[      84] = 32'h0;  // 32'hb0771b4c;
    ram_cell[      85] = 32'h0;  // 32'h5e64ccf8;
    ram_cell[      86] = 32'h0;  // 32'h08007872;
    ram_cell[      87] = 32'h0;  // 32'hb815abb2;
    ram_cell[      88] = 32'h0;  // 32'ha7b5e602;
    ram_cell[      89] = 32'h0;  // 32'he04d51e7;
    ram_cell[      90] = 32'h0;  // 32'h0db19ecd;
    ram_cell[      91] = 32'h0;  // 32'h18fc65bd;
    ram_cell[      92] = 32'h0;  // 32'h6560f8b8;
    ram_cell[      93] = 32'h0;  // 32'hcfed1dd6;
    ram_cell[      94] = 32'h0;  // 32'h2765c771;
    ram_cell[      95] = 32'h0;  // 32'h7459b8a5;
    ram_cell[      96] = 32'h0;  // 32'he45e6202;
    ram_cell[      97] = 32'h0;  // 32'hce758800;
    ram_cell[      98] = 32'h0;  // 32'h8dbac278;
    ram_cell[      99] = 32'h0;  // 32'h295bbabc;
    ram_cell[     100] = 32'h0;  // 32'h89ad71bc;
    ram_cell[     101] = 32'h0;  // 32'h1064ce51;
    ram_cell[     102] = 32'h0;  // 32'h477502a9;
    ram_cell[     103] = 32'h0;  // 32'h63ac3258;
    ram_cell[     104] = 32'h0;  // 32'h58ce5053;
    ram_cell[     105] = 32'h0;  // 32'h6d9ad95e;
    ram_cell[     106] = 32'h0;  // 32'hbcd7baa9;
    ram_cell[     107] = 32'h0;  // 32'hb69bdaef;
    ram_cell[     108] = 32'h0;  // 32'h990c2ff1;
    ram_cell[     109] = 32'h0;  // 32'h4e49e898;
    ram_cell[     110] = 32'h0;  // 32'h3ad49159;
    ram_cell[     111] = 32'h0;  // 32'h121fe1fa;
    ram_cell[     112] = 32'h0;  // 32'hcf5ed4aa;
    ram_cell[     113] = 32'h0;  // 32'h03151a71;
    ram_cell[     114] = 32'h0;  // 32'hd753a989;
    ram_cell[     115] = 32'h0;  // 32'h9756c828;
    ram_cell[     116] = 32'h0;  // 32'h39893111;
    ram_cell[     117] = 32'h0;  // 32'h14c678fa;
    ram_cell[     118] = 32'h0;  // 32'h15e90795;
    ram_cell[     119] = 32'h0;  // 32'h45076e70;
    ram_cell[     120] = 32'h0;  // 32'h4b38bc1e;
    ram_cell[     121] = 32'h0;  // 32'he7a5fd02;
    ram_cell[     122] = 32'h0;  // 32'h5925c265;
    ram_cell[     123] = 32'h0;  // 32'h19baa0cd;
    ram_cell[     124] = 32'h0;  // 32'h43f57f3a;
    ram_cell[     125] = 32'h0;  // 32'h0fed1ea1;
    ram_cell[     126] = 32'h0;  // 32'h497febe8;
    ram_cell[     127] = 32'h0;  // 32'h9218d3bf;
    ram_cell[     128] = 32'h0;  // 32'h01e2b55c;
    ram_cell[     129] = 32'h0;  // 32'hbc4d09a2;
    ram_cell[     130] = 32'h0;  // 32'h91e1392b;
    ram_cell[     131] = 32'h0;  // 32'h63c73d30;
    ram_cell[     132] = 32'h0;  // 32'hc0a0a0e6;
    ram_cell[     133] = 32'h0;  // 32'hea8ee38d;
    ram_cell[     134] = 32'h0;  // 32'h33d6b167;
    ram_cell[     135] = 32'h0;  // 32'h54ad4152;
    ram_cell[     136] = 32'h0;  // 32'hc9e9e92f;
    ram_cell[     137] = 32'h0;  // 32'h32579122;
    ram_cell[     138] = 32'h0;  // 32'h8f9e0e71;
    ram_cell[     139] = 32'h0;  // 32'h049e065b;
    ram_cell[     140] = 32'h0;  // 32'h170f3568;
    ram_cell[     141] = 32'h0;  // 32'hed2dc1bb;
    ram_cell[     142] = 32'h0;  // 32'h93df1b53;
    ram_cell[     143] = 32'h0;  // 32'ha1da44a3;
    ram_cell[     144] = 32'h0;  // 32'had9463e7;
    ram_cell[     145] = 32'h0;  // 32'haaabe717;
    ram_cell[     146] = 32'h0;  // 32'ha4e2e4c3;
    ram_cell[     147] = 32'h0;  // 32'h4b65b2f9;
    ram_cell[     148] = 32'h0;  // 32'he0cbcca3;
    ram_cell[     149] = 32'h0;  // 32'hac9fb9d3;
    ram_cell[     150] = 32'h0;  // 32'hf95101f7;
    ram_cell[     151] = 32'h0;  // 32'h6f59590c;
    ram_cell[     152] = 32'h0;  // 32'h13761f2b;
    ram_cell[     153] = 32'h0;  // 32'h219f6c2a;
    ram_cell[     154] = 32'h0;  // 32'h322e9677;
    ram_cell[     155] = 32'h0;  // 32'hb1f5c936;
    ram_cell[     156] = 32'h0;  // 32'hb0caa05b;
    ram_cell[     157] = 32'h0;  // 32'he370eb6b;
    ram_cell[     158] = 32'h0;  // 32'ha9d39ad6;
    ram_cell[     159] = 32'h0;  // 32'hbceaf300;
    ram_cell[     160] = 32'h0;  // 32'ha13ad4b5;
    ram_cell[     161] = 32'h0;  // 32'h33bbc9f0;
    ram_cell[     162] = 32'h0;  // 32'h562464f2;
    ram_cell[     163] = 32'h0;  // 32'hdfeafd8e;
    ram_cell[     164] = 32'h0;  // 32'h680e7a8d;
    ram_cell[     165] = 32'h0;  // 32'hfbf270d5;
    ram_cell[     166] = 32'h0;  // 32'h8eb70ecd;
    ram_cell[     167] = 32'h0;  // 32'h24f07199;
    ram_cell[     168] = 32'h0;  // 32'h9784c205;
    ram_cell[     169] = 32'h0;  // 32'h911d3f5a;
    ram_cell[     170] = 32'h0;  // 32'heea4d562;
    ram_cell[     171] = 32'h0;  // 32'h5b05e25f;
    ram_cell[     172] = 32'h0;  // 32'h94d6084b;
    ram_cell[     173] = 32'h0;  // 32'h019c96d1;
    ram_cell[     174] = 32'h0;  // 32'hf8c09bfd;
    ram_cell[     175] = 32'h0;  // 32'hc1aa4327;
    ram_cell[     176] = 32'h0;  // 32'hee0cfb91;
    ram_cell[     177] = 32'h0;  // 32'he4828172;
    ram_cell[     178] = 32'h0;  // 32'hd379e5e8;
    ram_cell[     179] = 32'h0;  // 32'h1d6e3c12;
    ram_cell[     180] = 32'h0;  // 32'h64c62186;
    ram_cell[     181] = 32'h0;  // 32'h8b8fe6ef;
    ram_cell[     182] = 32'h0;  // 32'hca9bb5af;
    ram_cell[     183] = 32'h0;  // 32'h9e5cc664;
    ram_cell[     184] = 32'h0;  // 32'h4bae7d16;
    ram_cell[     185] = 32'h0;  // 32'habb562a8;
    ram_cell[     186] = 32'h0;  // 32'hfc885cbb;
    ram_cell[     187] = 32'h0;  // 32'hd05e90ad;
    ram_cell[     188] = 32'h0;  // 32'h3d58fb38;
    ram_cell[     189] = 32'h0;  // 32'haed90805;
    ram_cell[     190] = 32'h0;  // 32'h276bd823;
    ram_cell[     191] = 32'h0;  // 32'h5ac35d38;
    ram_cell[     192] = 32'h0;  // 32'h2190ac74;
    ram_cell[     193] = 32'h0;  // 32'h793bd63e;
    ram_cell[     194] = 32'h0;  // 32'h1da46429;
    ram_cell[     195] = 32'h0;  // 32'h59daba02;
    ram_cell[     196] = 32'h0;  // 32'h41f9ccbf;
    ram_cell[     197] = 32'h0;  // 32'h89cc95ba;
    ram_cell[     198] = 32'h0;  // 32'h2f103508;
    ram_cell[     199] = 32'h0;  // 32'h0b3625a4;
    ram_cell[     200] = 32'h0;  // 32'he82d6218;
    ram_cell[     201] = 32'h0;  // 32'hf4211023;
    ram_cell[     202] = 32'h0;  // 32'h2a7973d2;
    ram_cell[     203] = 32'h0;  // 32'h2eb1e4d8;
    ram_cell[     204] = 32'h0;  // 32'h339768cd;
    ram_cell[     205] = 32'h0;  // 32'hc649ed0d;
    ram_cell[     206] = 32'h0;  // 32'h277e9475;
    ram_cell[     207] = 32'h0;  // 32'h2d92300e;
    ram_cell[     208] = 32'h0;  // 32'h0f9e4355;
    ram_cell[     209] = 32'h0;  // 32'hfc0c2482;
    ram_cell[     210] = 32'h0;  // 32'h09670c03;
    ram_cell[     211] = 32'h0;  // 32'h3120768c;
    ram_cell[     212] = 32'h0;  // 32'h80a86d37;
    ram_cell[     213] = 32'h0;  // 32'hbf414ec1;
    ram_cell[     214] = 32'h0;  // 32'hdf825577;
    ram_cell[     215] = 32'h0;  // 32'hea93f63a;
    ram_cell[     216] = 32'h0;  // 32'h3c4d124c;
    ram_cell[     217] = 32'h0;  // 32'h32cabbd3;
    ram_cell[     218] = 32'h0;  // 32'hdca3575f;
    ram_cell[     219] = 32'h0;  // 32'hb078ecc3;
    ram_cell[     220] = 32'h0;  // 32'h283a88af;
    ram_cell[     221] = 32'h0;  // 32'hafc3fa95;
    ram_cell[     222] = 32'h0;  // 32'he5d1f266;
    ram_cell[     223] = 32'h0;  // 32'h6dde6035;
    ram_cell[     224] = 32'h0;  // 32'hc0876400;
    ram_cell[     225] = 32'h0;  // 32'h46b7ff6f;
    ram_cell[     226] = 32'h0;  // 32'hdc5c2cb2;
    ram_cell[     227] = 32'h0;  // 32'hf1ceebcc;
    ram_cell[     228] = 32'h0;  // 32'h907c34a3;
    ram_cell[     229] = 32'h0;  // 32'h52322382;
    ram_cell[     230] = 32'h0;  // 32'hb99daa77;
    ram_cell[     231] = 32'h0;  // 32'h5aaad9ff;
    ram_cell[     232] = 32'h0;  // 32'h4e056a0e;
    ram_cell[     233] = 32'h0;  // 32'hb712c11f;
    ram_cell[     234] = 32'h0;  // 32'h18873c81;
    ram_cell[     235] = 32'h0;  // 32'haafe0593;
    ram_cell[     236] = 32'h0;  // 32'h0d2dc2d5;
    ram_cell[     237] = 32'h0;  // 32'h77259a84;
    ram_cell[     238] = 32'h0;  // 32'hd68e97ca;
    ram_cell[     239] = 32'h0;  // 32'h26988862;
    ram_cell[     240] = 32'h0;  // 32'he0ee5ee1;
    ram_cell[     241] = 32'h0;  // 32'h57037384;
    ram_cell[     242] = 32'h0;  // 32'hfa63129c;
    ram_cell[     243] = 32'h0;  // 32'h57e53da5;
    ram_cell[     244] = 32'h0;  // 32'hb4f74340;
    ram_cell[     245] = 32'h0;  // 32'h5a465b8d;
    ram_cell[     246] = 32'h0;  // 32'hb8c7102a;
    ram_cell[     247] = 32'h0;  // 32'hbd13d05a;
    ram_cell[     248] = 32'h0;  // 32'h26042a53;
    ram_cell[     249] = 32'h0;  // 32'h54ad1028;
    ram_cell[     250] = 32'h0;  // 32'h0a2533e3;
    ram_cell[     251] = 32'h0;  // 32'h64a52e62;
    ram_cell[     252] = 32'h0;  // 32'ha9f5ac5c;
    ram_cell[     253] = 32'h0;  // 32'he9a179a8;
    ram_cell[     254] = 32'h0;  // 32'h9a57aa1e;
    ram_cell[     255] = 32'h0;  // 32'h1324b5ec;
    // src matrix A
    ram_cell[     256] = 32'h2c6b1c5d;
    ram_cell[     257] = 32'ha513af34;
    ram_cell[     258] = 32'h0062a322;
    ram_cell[     259] = 32'h778b1a77;
    ram_cell[     260] = 32'heb95c33c;
    ram_cell[     261] = 32'hb73ffba4;
    ram_cell[     262] = 32'h771526be;
    ram_cell[     263] = 32'h910bc430;
    ram_cell[     264] = 32'hf6d71ed4;
    ram_cell[     265] = 32'h02f3ad4d;
    ram_cell[     266] = 32'h2254392a;
    ram_cell[     267] = 32'ha5780ef2;
    ram_cell[     268] = 32'hce810f6f;
    ram_cell[     269] = 32'h0f92cf0d;
    ram_cell[     270] = 32'h2330a974;
    ram_cell[     271] = 32'hce2893eb;
    ram_cell[     272] = 32'h1754e0fa;
    ram_cell[     273] = 32'hfa57d871;
    ram_cell[     274] = 32'heb59c353;
    ram_cell[     275] = 32'h72fad79b;
    ram_cell[     276] = 32'hc4ec54e5;
    ram_cell[     277] = 32'h2bfc5b3e;
    ram_cell[     278] = 32'h744a6453;
    ram_cell[     279] = 32'hffc79b0e;
    ram_cell[     280] = 32'h02d1ccd7;
    ram_cell[     281] = 32'h362dc9df;
    ram_cell[     282] = 32'hebc7529d;
    ram_cell[     283] = 32'ha8e3c9df;
    ram_cell[     284] = 32'h58fb37f5;
    ram_cell[     285] = 32'h2905b340;
    ram_cell[     286] = 32'he32a1441;
    ram_cell[     287] = 32'h178c67a6;
    ram_cell[     288] = 32'he36d9b71;
    ram_cell[     289] = 32'hb121628e;
    ram_cell[     290] = 32'hc7bfc646;
    ram_cell[     291] = 32'h640ae20f;
    ram_cell[     292] = 32'h500faa70;
    ram_cell[     293] = 32'ha7713970;
    ram_cell[     294] = 32'h1a2e93f3;
    ram_cell[     295] = 32'h4e035c7c;
    ram_cell[     296] = 32'h3a36048c;
    ram_cell[     297] = 32'h4e7b62ed;
    ram_cell[     298] = 32'h475d13a5;
    ram_cell[     299] = 32'he23a92cc;
    ram_cell[     300] = 32'h64203139;
    ram_cell[     301] = 32'ha0697ff9;
    ram_cell[     302] = 32'ha2d3433f;
    ram_cell[     303] = 32'hdb933dfd;
    ram_cell[     304] = 32'h6eb802bf;
    ram_cell[     305] = 32'hb9fe4c7b;
    ram_cell[     306] = 32'hd9e37223;
    ram_cell[     307] = 32'h4537a1ef;
    ram_cell[     308] = 32'h1d6b69c4;
    ram_cell[     309] = 32'hda317c7a;
    ram_cell[     310] = 32'h88617616;
    ram_cell[     311] = 32'h6030b3d7;
    ram_cell[     312] = 32'ha23b48c2;
    ram_cell[     313] = 32'h15bbbb8a;
    ram_cell[     314] = 32'h9ec2f717;
    ram_cell[     315] = 32'h79f39655;
    ram_cell[     316] = 32'h8af3ad4e;
    ram_cell[     317] = 32'h8c6c796c;
    ram_cell[     318] = 32'h0d16e125;
    ram_cell[     319] = 32'h4968efd1;
    ram_cell[     320] = 32'h22b877a3;
    ram_cell[     321] = 32'h67245a11;
    ram_cell[     322] = 32'hc815fb03;
    ram_cell[     323] = 32'hb1308acb;
    ram_cell[     324] = 32'h19fb6cbd;
    ram_cell[     325] = 32'h3d4fd17c;
    ram_cell[     326] = 32'h82144d63;
    ram_cell[     327] = 32'ha677284e;
    ram_cell[     328] = 32'h2a6310e7;
    ram_cell[     329] = 32'h0e6395b6;
    ram_cell[     330] = 32'hc754721b;
    ram_cell[     331] = 32'h0c943a5e;
    ram_cell[     332] = 32'h11be170d;
    ram_cell[     333] = 32'ha686eb5a;
    ram_cell[     334] = 32'h2805aa9e;
    ram_cell[     335] = 32'ha31abece;
    ram_cell[     336] = 32'he8235ee0;
    ram_cell[     337] = 32'hb4c64a2c;
    ram_cell[     338] = 32'h47c7f412;
    ram_cell[     339] = 32'h1d19ed11;
    ram_cell[     340] = 32'haa9d8d3e;
    ram_cell[     341] = 32'hb999b65b;
    ram_cell[     342] = 32'h24669007;
    ram_cell[     343] = 32'hbf067fb0;
    ram_cell[     344] = 32'h610b88d2;
    ram_cell[     345] = 32'h1bfb02fa;
    ram_cell[     346] = 32'hee754416;
    ram_cell[     347] = 32'h07c78f65;
    ram_cell[     348] = 32'h56aaa362;
    ram_cell[     349] = 32'h2981b3f3;
    ram_cell[     350] = 32'h328afd97;
    ram_cell[     351] = 32'h60fe2997;
    ram_cell[     352] = 32'hf05c0f99;
    ram_cell[     353] = 32'hb3bf7e73;
    ram_cell[     354] = 32'h5652431e;
    ram_cell[     355] = 32'he3c5725c;
    ram_cell[     356] = 32'hb5db8f78;
    ram_cell[     357] = 32'h2e13fdf3;
    ram_cell[     358] = 32'h0fe5ea0a;
    ram_cell[     359] = 32'hd4c3e5ae;
    ram_cell[     360] = 32'hdeb55f63;
    ram_cell[     361] = 32'h6b8b40f9;
    ram_cell[     362] = 32'h3721ce69;
    ram_cell[     363] = 32'h5b5b6761;
    ram_cell[     364] = 32'hda34cddb;
    ram_cell[     365] = 32'h8798daca;
    ram_cell[     366] = 32'hf9f6f878;
    ram_cell[     367] = 32'h84ad5748;
    ram_cell[     368] = 32'h80774ecd;
    ram_cell[     369] = 32'hdadfbe3a;
    ram_cell[     370] = 32'h40efc125;
    ram_cell[     371] = 32'h348f8a8f;
    ram_cell[     372] = 32'hbae5dc8d;
    ram_cell[     373] = 32'hdb1ae093;
    ram_cell[     374] = 32'h2d18654d;
    ram_cell[     375] = 32'h17625749;
    ram_cell[     376] = 32'h86bc909f;
    ram_cell[     377] = 32'h191f858c;
    ram_cell[     378] = 32'h9c28fc37;
    ram_cell[     379] = 32'hebdb5daf;
    ram_cell[     380] = 32'h15cf0197;
    ram_cell[     381] = 32'h63091964;
    ram_cell[     382] = 32'h74b9d837;
    ram_cell[     383] = 32'h20404647;
    ram_cell[     384] = 32'hd7af3fd4;
    ram_cell[     385] = 32'h3a4933f2;
    ram_cell[     386] = 32'h7b5eee7e;
    ram_cell[     387] = 32'haafa602b;
    ram_cell[     388] = 32'h4f8d3ee6;
    ram_cell[     389] = 32'h711cc234;
    ram_cell[     390] = 32'h9bfec07c;
    ram_cell[     391] = 32'h5694f6a3;
    ram_cell[     392] = 32'h65663661;
    ram_cell[     393] = 32'h908a32d0;
    ram_cell[     394] = 32'hc44c59b8;
    ram_cell[     395] = 32'h19e8bd7c;
    ram_cell[     396] = 32'h68c17606;
    ram_cell[     397] = 32'hd5fc22b3;
    ram_cell[     398] = 32'ha46f9bf3;
    ram_cell[     399] = 32'h3fcb7502;
    ram_cell[     400] = 32'hf2e51238;
    ram_cell[     401] = 32'he9955027;
    ram_cell[     402] = 32'hb62d9c14;
    ram_cell[     403] = 32'h2c81f127;
    ram_cell[     404] = 32'hbde894a8;
    ram_cell[     405] = 32'h307f4598;
    ram_cell[     406] = 32'h6e381e2e;
    ram_cell[     407] = 32'h7c1ffe04;
    ram_cell[     408] = 32'he52fe1a9;
    ram_cell[     409] = 32'he25f4077;
    ram_cell[     410] = 32'h3327e419;
    ram_cell[     411] = 32'hb3108b91;
    ram_cell[     412] = 32'h96834c89;
    ram_cell[     413] = 32'h72be8954;
    ram_cell[     414] = 32'h17891cb2;
    ram_cell[     415] = 32'h5487fa44;
    ram_cell[     416] = 32'h8aa533a0;
    ram_cell[     417] = 32'hc1ed6f94;
    ram_cell[     418] = 32'h0ad3e50e;
    ram_cell[     419] = 32'he1d9194b;
    ram_cell[     420] = 32'hb12718f8;
    ram_cell[     421] = 32'h430fed16;
    ram_cell[     422] = 32'h5b61d106;
    ram_cell[     423] = 32'h352e0b8a;
    ram_cell[     424] = 32'hb3573abb;
    ram_cell[     425] = 32'hf94a6529;
    ram_cell[     426] = 32'hca898aeb;
    ram_cell[     427] = 32'h3960cd4d;
    ram_cell[     428] = 32'hcd110ae5;
    ram_cell[     429] = 32'hc650831b;
    ram_cell[     430] = 32'h5e59a2b7;
    ram_cell[     431] = 32'ha2cee168;
    ram_cell[     432] = 32'hc969cb13;
    ram_cell[     433] = 32'hff44d0ce;
    ram_cell[     434] = 32'hb8714d05;
    ram_cell[     435] = 32'h3bc0f871;
    ram_cell[     436] = 32'hb94ff94b;
    ram_cell[     437] = 32'h7cf95d45;
    ram_cell[     438] = 32'h5e95d197;
    ram_cell[     439] = 32'h79a702d0;
    ram_cell[     440] = 32'hed182597;
    ram_cell[     441] = 32'h061617f7;
    ram_cell[     442] = 32'had3af8c2;
    ram_cell[     443] = 32'h37504a07;
    ram_cell[     444] = 32'ha5830c11;
    ram_cell[     445] = 32'hcf6025e5;
    ram_cell[     446] = 32'h385ae034;
    ram_cell[     447] = 32'h8617697d;
    ram_cell[     448] = 32'h4e0556d9;
    ram_cell[     449] = 32'ha4e98324;
    ram_cell[     450] = 32'h30c3ed19;
    ram_cell[     451] = 32'hb951535a;
    ram_cell[     452] = 32'hf2766c8e;
    ram_cell[     453] = 32'h3fa6434a;
    ram_cell[     454] = 32'hce56c887;
    ram_cell[     455] = 32'h35a9f898;
    ram_cell[     456] = 32'hcde30561;
    ram_cell[     457] = 32'hc15467c9;
    ram_cell[     458] = 32'h0d4224fc;
    ram_cell[     459] = 32'hd7f4dd7d;
    ram_cell[     460] = 32'h9368da22;
    ram_cell[     461] = 32'hbaecf542;
    ram_cell[     462] = 32'h518e019a;
    ram_cell[     463] = 32'h34e18386;
    ram_cell[     464] = 32'hb5629917;
    ram_cell[     465] = 32'h39da3d20;
    ram_cell[     466] = 32'h485d5606;
    ram_cell[     467] = 32'h5ad56b48;
    ram_cell[     468] = 32'he0e0070f;
    ram_cell[     469] = 32'h075ef9b7;
    ram_cell[     470] = 32'h2c47d4db;
    ram_cell[     471] = 32'hfa0edaac;
    ram_cell[     472] = 32'h5fc12578;
    ram_cell[     473] = 32'hdb23b8cb;
    ram_cell[     474] = 32'hf53ea79d;
    ram_cell[     475] = 32'h357dea6b;
    ram_cell[     476] = 32'h3d105ef2;
    ram_cell[     477] = 32'h328fd3c2;
    ram_cell[     478] = 32'hf6ab7608;
    ram_cell[     479] = 32'h472741fe;
    ram_cell[     480] = 32'h2321228d;
    ram_cell[     481] = 32'h5f065b42;
    ram_cell[     482] = 32'he048e334;
    ram_cell[     483] = 32'h36f55c7e;
    ram_cell[     484] = 32'hbcda1a84;
    ram_cell[     485] = 32'hea602362;
    ram_cell[     486] = 32'h61ea4052;
    ram_cell[     487] = 32'h88cbc117;
    ram_cell[     488] = 32'h8a167cd3;
    ram_cell[     489] = 32'hff999006;
    ram_cell[     490] = 32'h680153f6;
    ram_cell[     491] = 32'h20327de0;
    ram_cell[     492] = 32'h9f191ebf;
    ram_cell[     493] = 32'h361db764;
    ram_cell[     494] = 32'h70010a12;
    ram_cell[     495] = 32'hb39fe3f9;
    ram_cell[     496] = 32'h6b92acbc;
    ram_cell[     497] = 32'h9c08f30b;
    ram_cell[     498] = 32'hacb9fecc;
    ram_cell[     499] = 32'h3cf8d288;
    ram_cell[     500] = 32'h389985a7;
    ram_cell[     501] = 32'h6732aa75;
    ram_cell[     502] = 32'h7974d34c;
    ram_cell[     503] = 32'h624f75eb;
    ram_cell[     504] = 32'he3da0778;
    ram_cell[     505] = 32'h8f5b3c6d;
    ram_cell[     506] = 32'h7db6935d;
    ram_cell[     507] = 32'hefaefb2d;
    ram_cell[     508] = 32'hce89b9c7;
    ram_cell[     509] = 32'h24d36189;
    ram_cell[     510] = 32'h631fdc7c;
    ram_cell[     511] = 32'hd868c634;
    // src matrix B
    ram_cell[     512] = 32'hb41e9913;
    ram_cell[     513] = 32'h298b4524;
    ram_cell[     514] = 32'h006ebec8;
    ram_cell[     515] = 32'he7e1cf50;
    ram_cell[     516] = 32'hd0b4d8f5;
    ram_cell[     517] = 32'ha35e4be3;
    ram_cell[     518] = 32'he12220fb;
    ram_cell[     519] = 32'h868f4209;
    ram_cell[     520] = 32'h9719231a;
    ram_cell[     521] = 32'hb8f7b5c8;
    ram_cell[     522] = 32'hc2ee05b0;
    ram_cell[     523] = 32'h126437d0;
    ram_cell[     524] = 32'h01ea1295;
    ram_cell[     525] = 32'h4445a02d;
    ram_cell[     526] = 32'h54c6910a;
    ram_cell[     527] = 32'h354c7694;
    ram_cell[     528] = 32'h2a9c29ef;
    ram_cell[     529] = 32'hd770fd1e;
    ram_cell[     530] = 32'h3b45616d;
    ram_cell[     531] = 32'h58d647f3;
    ram_cell[     532] = 32'h00e20ef7;
    ram_cell[     533] = 32'hb6f332dd;
    ram_cell[     534] = 32'h09b9a645;
    ram_cell[     535] = 32'h9c43c594;
    ram_cell[     536] = 32'h66f3a33d;
    ram_cell[     537] = 32'heac152ca;
    ram_cell[     538] = 32'hfeaec8d0;
    ram_cell[     539] = 32'h16fb1ec8;
    ram_cell[     540] = 32'ha8af1760;
    ram_cell[     541] = 32'h94806cb9;
    ram_cell[     542] = 32'h5b3a5130;
    ram_cell[     543] = 32'hc92bb682;
    ram_cell[     544] = 32'hd3587a81;
    ram_cell[     545] = 32'h3cae7cf2;
    ram_cell[     546] = 32'hcfc0fa11;
    ram_cell[     547] = 32'h89094a60;
    ram_cell[     548] = 32'h7421f183;
    ram_cell[     549] = 32'h5375fd19;
    ram_cell[     550] = 32'hfe0b28ad;
    ram_cell[     551] = 32'h4d457c88;
    ram_cell[     552] = 32'h40d4ab0c;
    ram_cell[     553] = 32'h3c3aed2d;
    ram_cell[     554] = 32'h52bdd126;
    ram_cell[     555] = 32'hbc71bbb7;
    ram_cell[     556] = 32'he4f68102;
    ram_cell[     557] = 32'hb996d0d1;
    ram_cell[     558] = 32'h7a31c960;
    ram_cell[     559] = 32'h38762a08;
    ram_cell[     560] = 32'h19802914;
    ram_cell[     561] = 32'h970cb01a;
    ram_cell[     562] = 32'h5f83634b;
    ram_cell[     563] = 32'hef770aae;
    ram_cell[     564] = 32'h4ca5bbc9;
    ram_cell[     565] = 32'hb36fa4e6;
    ram_cell[     566] = 32'h2a79abd8;
    ram_cell[     567] = 32'h8852dee5;
    ram_cell[     568] = 32'ha8d94d14;
    ram_cell[     569] = 32'he9e492ee;
    ram_cell[     570] = 32'h7f6a0a0e;
    ram_cell[     571] = 32'hc10e4f4f;
    ram_cell[     572] = 32'hc8138d39;
    ram_cell[     573] = 32'h1d53915d;
    ram_cell[     574] = 32'h5645307d;
    ram_cell[     575] = 32'hf228f462;
    ram_cell[     576] = 32'h4dcc01c7;
    ram_cell[     577] = 32'hff8814c4;
    ram_cell[     578] = 32'h03ec58b4;
    ram_cell[     579] = 32'h89f33f2e;
    ram_cell[     580] = 32'hebbf6fb0;
    ram_cell[     581] = 32'hcbd8994b;
    ram_cell[     582] = 32'hbd1f174f;
    ram_cell[     583] = 32'hbdfc7b23;
    ram_cell[     584] = 32'h55b559ba;
    ram_cell[     585] = 32'hfe9be5bb;
    ram_cell[     586] = 32'h8372a549;
    ram_cell[     587] = 32'h05b112a9;
    ram_cell[     588] = 32'h0d1c52e1;
    ram_cell[     589] = 32'hd767b794;
    ram_cell[     590] = 32'h934535dc;
    ram_cell[     591] = 32'h33fa76c9;
    ram_cell[     592] = 32'hb5b5c504;
    ram_cell[     593] = 32'h0e08177f;
    ram_cell[     594] = 32'h96af52f0;
    ram_cell[     595] = 32'h324ee929;
    ram_cell[     596] = 32'hda4820a1;
    ram_cell[     597] = 32'h10c2b407;
    ram_cell[     598] = 32'h89549e2d;
    ram_cell[     599] = 32'h038a5f3a;
    ram_cell[     600] = 32'h97490256;
    ram_cell[     601] = 32'hc5710b6c;
    ram_cell[     602] = 32'h83ee5e28;
    ram_cell[     603] = 32'hc77b94dc;
    ram_cell[     604] = 32'h9a08ee30;
    ram_cell[     605] = 32'hed6419e9;
    ram_cell[     606] = 32'h8f08c106;
    ram_cell[     607] = 32'h865b222e;
    ram_cell[     608] = 32'hf9a7e585;
    ram_cell[     609] = 32'h13a43193;
    ram_cell[     610] = 32'h7245bf97;
    ram_cell[     611] = 32'h48d002a9;
    ram_cell[     612] = 32'h523a500e;
    ram_cell[     613] = 32'hbe145629;
    ram_cell[     614] = 32'h63a742d9;
    ram_cell[     615] = 32'h1c97e1de;
    ram_cell[     616] = 32'hb0cf89c0;
    ram_cell[     617] = 32'hc6685f6e;
    ram_cell[     618] = 32'h2bdf1475;
    ram_cell[     619] = 32'hcb14c1b2;
    ram_cell[     620] = 32'he056fcf9;
    ram_cell[     621] = 32'hec1e03ae;
    ram_cell[     622] = 32'h34286cb4;
    ram_cell[     623] = 32'hd2671c38;
    ram_cell[     624] = 32'h48eadd14;
    ram_cell[     625] = 32'h9ac4ebb4;
    ram_cell[     626] = 32'h6e077961;
    ram_cell[     627] = 32'hd3c79255;
    ram_cell[     628] = 32'h326a2231;
    ram_cell[     629] = 32'h9d74f67b;
    ram_cell[     630] = 32'hc24064f3;
    ram_cell[     631] = 32'hffcf328d;
    ram_cell[     632] = 32'he970c466;
    ram_cell[     633] = 32'h25ce163e;
    ram_cell[     634] = 32'h3bbb3a12;
    ram_cell[     635] = 32'he78fe247;
    ram_cell[     636] = 32'h52eaa932;
    ram_cell[     637] = 32'h4f434e7d;
    ram_cell[     638] = 32'h391c4c5f;
    ram_cell[     639] = 32'he0d975a9;
    ram_cell[     640] = 32'h13255069;
    ram_cell[     641] = 32'hb9c8a357;
    ram_cell[     642] = 32'h76fab913;
    ram_cell[     643] = 32'h5c5f841b;
    ram_cell[     644] = 32'hf8fbe619;
    ram_cell[     645] = 32'h3c1ea5b7;
    ram_cell[     646] = 32'h98714baf;
    ram_cell[     647] = 32'h5ec02ffd;
    ram_cell[     648] = 32'hc1c52548;
    ram_cell[     649] = 32'hf883c676;
    ram_cell[     650] = 32'h6648cd62;
    ram_cell[     651] = 32'h73672094;
    ram_cell[     652] = 32'h7f9df761;
    ram_cell[     653] = 32'h3687e5f8;
    ram_cell[     654] = 32'h21fe6cde;
    ram_cell[     655] = 32'h64f75fc5;
    ram_cell[     656] = 32'hde764fb0;
    ram_cell[     657] = 32'hf108e500;
    ram_cell[     658] = 32'h3a98426e;
    ram_cell[     659] = 32'h5a7c8855;
    ram_cell[     660] = 32'h5a0924fe;
    ram_cell[     661] = 32'h2bc650ee;
    ram_cell[     662] = 32'he41eae9b;
    ram_cell[     663] = 32'h5aee70d8;
    ram_cell[     664] = 32'h0476be11;
    ram_cell[     665] = 32'ha0adad9a;
    ram_cell[     666] = 32'h4acb72b9;
    ram_cell[     667] = 32'hcecf1597;
    ram_cell[     668] = 32'he779f9de;
    ram_cell[     669] = 32'h70e86f2a;
    ram_cell[     670] = 32'h005863f0;
    ram_cell[     671] = 32'h3e9cc738;
    ram_cell[     672] = 32'hec44e2f6;
    ram_cell[     673] = 32'h390e027c;
    ram_cell[     674] = 32'h5fdd73b8;
    ram_cell[     675] = 32'h171e13b4;
    ram_cell[     676] = 32'h0fc59d91;
    ram_cell[     677] = 32'hae1abee5;
    ram_cell[     678] = 32'h6a7325b1;
    ram_cell[     679] = 32'h48245ece;
    ram_cell[     680] = 32'h5fbb3c66;
    ram_cell[     681] = 32'h1f4ac2cc;
    ram_cell[     682] = 32'h96ef2408;
    ram_cell[     683] = 32'h05a973b7;
    ram_cell[     684] = 32'h0b53e838;
    ram_cell[     685] = 32'hb13ba0ea;
    ram_cell[     686] = 32'h9bb32a19;
    ram_cell[     687] = 32'h69cddff1;
    ram_cell[     688] = 32'h12f0d512;
    ram_cell[     689] = 32'hc915ca8c;
    ram_cell[     690] = 32'hf9cc9036;
    ram_cell[     691] = 32'h34390071;
    ram_cell[     692] = 32'hf5ae7ee0;
    ram_cell[     693] = 32'hb84052ec;
    ram_cell[     694] = 32'ha8847cd7;
    ram_cell[     695] = 32'ha3fc51ca;
    ram_cell[     696] = 32'h42bb72db;
    ram_cell[     697] = 32'hf711535a;
    ram_cell[     698] = 32'h062e658c;
    ram_cell[     699] = 32'h5fc4c91c;
    ram_cell[     700] = 32'hfeb2776c;
    ram_cell[     701] = 32'h8d56f2f3;
    ram_cell[     702] = 32'h8b83a52d;
    ram_cell[     703] = 32'hfabd87b1;
    ram_cell[     704] = 32'h0d60b66f;
    ram_cell[     705] = 32'h42892270;
    ram_cell[     706] = 32'h5899e40e;
    ram_cell[     707] = 32'h591ca4a3;
    ram_cell[     708] = 32'hf8ed9fbd;
    ram_cell[     709] = 32'h73cf3830;
    ram_cell[     710] = 32'h0e820666;
    ram_cell[     711] = 32'ha27dcc7e;
    ram_cell[     712] = 32'h50d18db0;
    ram_cell[     713] = 32'hc6b92b98;
    ram_cell[     714] = 32'h51b47b4e;
    ram_cell[     715] = 32'ha2e1ba9f;
    ram_cell[     716] = 32'h3c208fe5;
    ram_cell[     717] = 32'hc4fd0c08;
    ram_cell[     718] = 32'h51e15205;
    ram_cell[     719] = 32'h990ce639;
    ram_cell[     720] = 32'hd6f68d0a;
    ram_cell[     721] = 32'he54771cd;
    ram_cell[     722] = 32'h5b8762c0;
    ram_cell[     723] = 32'hc6532bdd;
    ram_cell[     724] = 32'hadc7143d;
    ram_cell[     725] = 32'had90569a;
    ram_cell[     726] = 32'hc3ed3959;
    ram_cell[     727] = 32'h12300bf4;
    ram_cell[     728] = 32'h9d3fbe50;
    ram_cell[     729] = 32'hae6fb823;
    ram_cell[     730] = 32'h36d96bbd;
    ram_cell[     731] = 32'h6f023425;
    ram_cell[     732] = 32'hdfd2ffa2;
    ram_cell[     733] = 32'h33b44f6e;
    ram_cell[     734] = 32'h0ed7d080;
    ram_cell[     735] = 32'hef666697;
    ram_cell[     736] = 32'h28616cef;
    ram_cell[     737] = 32'hf30f6060;
    ram_cell[     738] = 32'h37089d3a;
    ram_cell[     739] = 32'haa6bc1fd;
    ram_cell[     740] = 32'h0fed7130;
    ram_cell[     741] = 32'hc3bd49bd;
    ram_cell[     742] = 32'hba0a5ff0;
    ram_cell[     743] = 32'hc1243eb5;
    ram_cell[     744] = 32'hfac8e0f9;
    ram_cell[     745] = 32'hb1ae530b;
    ram_cell[     746] = 32'hf3459950;
    ram_cell[     747] = 32'hde650f28;
    ram_cell[     748] = 32'h57115822;
    ram_cell[     749] = 32'he749722d;
    ram_cell[     750] = 32'h99697bc3;
    ram_cell[     751] = 32'h6be516e8;
    ram_cell[     752] = 32'h2b4b7ea9;
    ram_cell[     753] = 32'h18b94a5e;
    ram_cell[     754] = 32'h44c09056;
    ram_cell[     755] = 32'ha66bf0e1;
    ram_cell[     756] = 32'hbe37b86b;
    ram_cell[     757] = 32'h8e80329b;
    ram_cell[     758] = 32'h7ed04642;
    ram_cell[     759] = 32'h5f4f8a16;
    ram_cell[     760] = 32'h43fe9e82;
    ram_cell[     761] = 32'h25351379;
    ram_cell[     762] = 32'h553a250d;
    ram_cell[     763] = 32'ha5c7bc69;
    ram_cell[     764] = 32'h957db63a;
    ram_cell[     765] = 32'h2d333e16;
    ram_cell[     766] = 32'h93ecbf74;
    ram_cell[     767] = 32'h5803133f;
end

endmodule

